--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A0000E0190001E0180001E0170003E0160005E015000AE0140013E0130020";
attribute INIT_01 of ram_1024_x_18  : label is "E9330900E9390900E937094DE010000E8001D0100113001AEE3D0E00EE3E0E00";
attribute INIT_02 of ram_1024_x_18  : label is "50314268623DEE3EAE00CE036E3EEE3D8E01CE036E3D0B130A080900E9350900";
attribute INIT_03 of ram_1024_x_18  : label is "404C50404401018B005A0100623D633EEF086F3EEF096F3D51994201623E4034";
attribute INIT_04 of ram_1024_x_18  : label is "00B40100623D633E4092CE086E08CE076E09EF086F3EEF096F3DC004E0240001";
attribute INIT_05 of ram_1024_x_18  : label is "CE076E09E009E108014A00B40100623D633EC004E0240002406350544401018B";
attribute INIT_06 of ram_1024_x_18  : label is "02B40300C004E0240003407A506B4401018B000E0101623D633E4092CE086E08";
attribute INIT_07 of ram_1024_x_18  : label is "613E020E0301C004E02400044092CE086E08CE076E09E009E108014A603D613E";
attribute INIT_08 of ram_1024_x_18  : label is "8F01EFFF6F08EF098F01EFFF6F094092CE086E08CE076E09E009E108014A603D";
attribute INIT_09 of ram_1024_x_18  : label is "50A3430013906139E1335498C301010A509B43001390613750D559A0A000EF08";
attribute INIT_0A of ram_1024_x_18  : label is "6039E037D0406435603750BB4480A4806408EF3B7F1011B0E13554A0C301010A";
attribute INIT_0B of ram_1024_x_18  : label is "6039E03790406435603740CAE108E009E100D020623B61086009E03990406433";
attribute INIT_0C of ram_1024_x_18  : label is "CE036E08CE036E098B018901E108E009A1009020623B61086009E039D0406433";
attribute INIT_0D of ram_1024_x_18  : label is "4003602440F4E0378001E0FF603740DE50D9400260244092C0066039C0056037";
attribute INIT_0E of ram_1024_x_18  : label is "603940F450EF4004602440F4E0398001E0FF6039E0378001E0FF603740EB50E2";
attribute INIT_0F of ram_1024_x_18  : label is "C002600BE0228028000A000AC001600DE00D6039E00B603740F4E0398001E0FF";
attribute INIT_10 of ram_1024_x_18  : label is "11601730162015101400401AC020003FC0176023C0166022E0238028000A000A";
attribute INIT_11 of ram_1024_x_18  : label is "10501170E004E105013710501160E002E103013710401170E000E10101371040";
attribute INIT_12 of ram_1024_x_18  : label is "6400650106000700018300006104620503000400650266030700E006E1070137";
attribute INIT_13 of ram_1024_x_18  : label is "931051403020040003000201E43DE33EE23FA000018304000500660667070183";
attribute INIT_14 of ram_1024_x_18  : label is "070014201530A000F130D020A000643D633E623F10401130553D020604080308";
attribute INIT_15 of ram_1024_x_18  : label is "56204177515F59755730A0004151A7008601F510D400595A5510E10054000600";
attribute INIT_16 of ram_1024_x_18  : label is "0804417D0801417D0802416F516B596D54004173516759715510417B51635979";
attribute INIT_17 of ram_1024_x_18  : label is "F150D040A000417D0804417D0801417D0804417D0801417D0804417D0801417D";
attribute INIT_18 of ram_1024_x_18  : label is "52004197518F59935310A000B1309020A000B370B260B1509040A000F370F260";
attribute INIT_19 of ram_1024_x_18  : label is "0000000000000000000000004199A00004044198040241980401419555975993";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "028E22B00A3DC0388AC028F700E22228F70088D3D2626008888A508888888888";
attribute INITP_01 of ram_1024_x_18 : label is "89A888E43D39090F4E43D388885A5024243A5024243420B6D0B6D0DA424388AC";
attribute INITP_02 of ram_1024_x_18 : label is "5B333333333F7F7F7F6D5754025800EA740AAC0300C0002B0AC2B0AC0038889A";
attribute INITP_03 of ram_1024_x_18 : label is "000000000000000000000000000000000000000000000000000E333F7F659565";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A0000E0190001E0180001E0170003E0160005E015000AE0140013E0130020",
                INIT_01 => X"E9330900E9390900E937094DE010000E8001D0100113001AEE3D0E00EE3E0E00",
                INIT_02 => X"50314268623DEE3EAE00CE036E3EEE3D8E01CE036E3D0B130A080900E9350900",
                INIT_03 => X"404C50404401018B005A0100623D633EEF086F3EEF096F3D51994201623E4034",
                INIT_04 => X"00B40100623D633E4092CE086E08CE076E09EF086F3EEF096F3DC004E0240001",
                INIT_05 => X"CE076E09E009E108014A00B40100623D633EC004E0240002406350544401018B",
                INIT_06 => X"02B40300C004E0240003407A506B4401018B000E0101623D633E4092CE086E08",
                INIT_07 => X"613E020E0301C004E02400044092CE086E08CE076E09E009E108014A603D613E",
                INIT_08 => X"8F01EFFF6F08EF098F01EFFF6F094092CE086E08CE076E09E009E108014A603D",
                INIT_09 => X"50A3430013906139E1335498C301010A509B43001390613750D559A0A000EF08",
                INIT_0A => X"6039E037D0406435603750BB4480A4806408EF3B7F1011B0E13554A0C301010A",
                INIT_0B => X"6039E03790406435603740CAE108E009E100D020623B61086009E03990406433",
                INIT_0C => X"CE036E08CE036E098B018901E108E009A1009020623B61086009E039D0406433",
                INIT_0D => X"4003602440F4E0378001E0FF603740DE50D9400260244092C0066039C0056037",
                INIT_0E => X"603940F450EF4004602440F4E0398001E0FF6039E0378001E0FF603740EB50E2",
                INIT_0F => X"C002600BE0228028000A000AC001600DE00D6039E00B603740F4E0398001E0FF",
                INIT_10 => X"11601730162015101400401AC020003FC0176023C0166022E0238028000A000A",
                INIT_11 => X"10501170E004E105013710501160E002E103013710401170E000E10101371040",
                INIT_12 => X"6400650106000700018300006104620503000400650266030700E006E1070137",
                INIT_13 => X"931051403020040003000201E43DE33EE23FA000018304000500660667070183",
                INIT_14 => X"070014201530A000F130D020A000643D633E623F10401130553D020604080308",
                INIT_15 => X"56204177515F59755730A0004151A7008601F510D400595A5510E10054000600",
                INIT_16 => X"0804417D0801417D0802416F516B596D54004173516759715510417B51635979",
                INIT_17 => X"F150D040A000417D0804417D0801417D0804417D0801417D0804417D0801417D",
                INIT_18 => X"52004197518F59935310A000B1309020A000B370B260B1509040A000F370F260",
                INIT_19 => X"0000000000000000000000004199A00004044198040241980401419555975993",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"028E22B00A3DC0388AC028F700E22228F70088D3D2626008888A508888888888",
               INITP_01 => X"89A888E43D39090F4E43D388885A5024243A5024243420B6D0B6D0DA424388AC",
               INITP_02 => X"5B333333333F7F7F7F6D5754025800EA740AAC0300C0002B0AC2B0AC0038889A",
               INITP_03 => X"000000000000000000000000000000000000000000000000000E333F7F659565",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
