--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E0190001E0180001E0170003E0160005E015000AE0140013E01300204001C001";
attribute INIT_01 of ram_1024_x_18  : label is "E9390900E937094DE010000E8001D0100113001AEE3D0E00EE3E0E00E01A0000";
attribute INIT_02 of ram_1024_x_18  : label is "EE3EAE00CE036E3EEE3D8E01C903CE036E3D0B130A080900E9350900E9330900";
attribute INIT_03 of ram_1024_x_18  : label is "018E005A0100623D633EEF086F3EEF096F3D519C4201623E403750344268623D";
attribute INIT_04 of ram_1024_x_18  : label is "633E4095CE086E08CE076E09EF086F3EEF096F3DC004E0240001404F50434401";
attribute INIT_05 of ram_1024_x_18  : label is "E108014D00B40100623D633EC004E0240002406650574401018E00B40100623D";
attribute INIT_06 of ram_1024_x_18  : label is "E0240003407D506E4401018E000E0101623D633E4095CE086E08CE076E09E009";
attribute INIT_07 of ram_1024_x_18  : label is "C004E02400044095CE086E08CE076E09E009E108014D603D613E02B40300C004";
attribute INIT_08 of ram_1024_x_18  : label is "EF098F01EFFF6F094095CE086E08CE076E09E009E108014D603D613E020E0301";
attribute INIT_09 of ram_1024_x_18  : label is "6139E133549BC301010A509E43001390613750D859A0A000EF088F01EFFF6F08";
attribute INIT_0A of ram_1024_x_18  : label is "6435603750BE4480A4806408EF3B7F1011B0E13554A3C301010A50A643001390";
attribute INIT_0B of ram_1024_x_18  : label is "6435603740CDE108E009E100D020623B61086009E039904064336039E037D040";
attribute INIT_0C of ram_1024_x_18  : label is "6E098B018901E108E009A1009020623B61086009E039D04064336039E0379040";
attribute INIT_0D of ram_1024_x_18  : label is "E0378001E0FF603740E150DC400260244095C0066039C0056037CE036E08CE03";
attribute INIT_0E of ram_1024_x_18  : label is "4004602440F7E0398001E0FF6039E0378001E0FF603740EE50E54003602440F7";
attribute INIT_0F of ram_1024_x_18  : label is "8028000A000AC001600DE00D6039E00B603740F7E0398001E0FF603940F750F2";
attribute INIT_10 of ram_1024_x_18  : label is "15101400401CC020003FC0176023C0166022E0238028000A000AC002600BE022";
attribute INIT_11 of ram_1024_x_18  : label is "E105013A10501160E002E103013A10401170E000E101013A1040116017301620";
attribute INIT_12 of ram_1024_x_18  : label is "0700018600006104620503000400650266030700E006E107013A10501170E004";
attribute INIT_13 of ram_1024_x_18  : label is "040003000201E43DE33EE23FA000018604000500660667070186640065010600";
attribute INIT_14 of ram_1024_x_18  : label is "A000F130D020A000643D633E623F104011305540020604080308931051433020";
attribute INIT_15 of ram_1024_x_18  : label is "59785730A0004154A7008601F510D400595D5510E10054000600070014201530";
attribute INIT_16 of ram_1024_x_18  : label is "418008024172516E597054004176516A59745510417E5166597C5620417A5162";
attribute INIT_17 of ram_1024_x_18  : label is "4180080441800801418008044180080141800804418008014180080441800801";
attribute INIT_18 of ram_1024_x_18  : label is "59965310A000B1309020A000B370B260B1509040A000F370F260F150D040A000";
attribute INIT_19 of ram_1024_x_18  : label is "4022C0164021419CA0000404419B0402419B04014198559A59965200419A5192";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000008001C020003FC017";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "419D000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "A388AC028F700E22B00A3DC038888A3DC02234F4989A008888A508888888888F";
attribute INITP_01 of ram_1024_x_18 : label is "6A22390F4E4243D390F4E222169409090E9409090D082DB42DB4369090E22B00";
attribute INITP_02 of ram_1024_x_18 : label is "CCCCCCCCCFDFDFDFDB55D50096003A9D02AB00C030000AC2B0AC2B000E2226A2";
attribute INITP_03 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000E2238CCFDFD9655956";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "C000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E0190001E0180001E0170003E0160005E015000AE0140013E01300204001C001",
                INIT_01 => X"E9390900E937094DE010000E8001D0100113001AEE3D0E00EE3E0E00E01A0000",
                INIT_02 => X"EE3EAE00CE036E3EEE3D8E01C903CE036E3D0B130A080900E9350900E9330900",
                INIT_03 => X"018E005A0100623D633EEF086F3EEF096F3D519C4201623E403750344268623D",
                INIT_04 => X"633E4095CE086E08CE076E09EF086F3EEF096F3DC004E0240001404F50434401",
                INIT_05 => X"E108014D00B40100623D633EC004E0240002406650574401018E00B40100623D",
                INIT_06 => X"E0240003407D506E4401018E000E0101623D633E4095CE086E08CE076E09E009",
                INIT_07 => X"C004E02400044095CE086E08CE076E09E009E108014D603D613E02B40300C004",
                INIT_08 => X"EF098F01EFFF6F094095CE086E08CE076E09E009E108014D603D613E020E0301",
                INIT_09 => X"6139E133549BC301010A509E43001390613750D859A0A000EF088F01EFFF6F08",
                INIT_0A => X"6435603750BE4480A4806408EF3B7F1011B0E13554A3C301010A50A643001390",
                INIT_0B => X"6435603740CDE108E009E100D020623B61086009E039904064336039E037D040",
                INIT_0C => X"6E098B018901E108E009A1009020623B61086009E039D04064336039E0379040",
                INIT_0D => X"E0378001E0FF603740E150DC400260244095C0066039C0056037CE036E08CE03",
                INIT_0E => X"4004602440F7E0398001E0FF6039E0378001E0FF603740EE50E54003602440F7",
                INIT_0F => X"8028000A000AC001600DE00D6039E00B603740F7E0398001E0FF603940F750F2",
                INIT_10 => X"15101400401CC020003FC0176023C0166022E0238028000A000AC002600BE022",
                INIT_11 => X"E105013A10501160E002E103013A10401170E000E101013A1040116017301620",
                INIT_12 => X"0700018600006104620503000400650266030700E006E107013A10501170E004",
                INIT_13 => X"040003000201E43DE33EE23FA000018604000500660667070186640065010600",
                INIT_14 => X"A000F130D020A000643D633E623F104011305540020604080308931051433020",
                INIT_15 => X"59785730A0004154A7008601F510D400595D5510E10054000600070014201530",
                INIT_16 => X"418008024172516E597054004176516A59745510417E5166597C5620417A5162",
                INIT_17 => X"4180080441800801418008044180080141800804418008014180080441800801",
                INIT_18 => X"59965310A000B1309020A000B370B260B1509040A000F370F260F150D040A000",
                INIT_19 => X"4022C0164021419CA0000404419B0402419B04014198559A59965200419A5192",
                INIT_1A => X"0000000000000000000000000000000000000000000000008001C020003FC017",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"419D000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"A388AC028F700E22B00A3DC038888A3DC02234F4989A008888A508888888888F",
               INITP_01 => X"6A22390F4E4243D390F4E222169409090E9409090D082DB42DB4369090E22B00",
               INITP_02 => X"CCCCCCCCCFDFDFDFDB55D50096003A9D02AB00C030000AC2B0AC2B000E2226A2",
               INITP_03 => X"0000000000000000000000000000000000000000000000E2238CCFDFD9655956",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"C000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
