--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A00D5E019001FE01800B6E017003EE01600B1E0150076E014000FE01300C9";
attribute INIT_01 of ram_1024_x_18  : label is "E02200FFE0210001E02000FFE01F0003E01E00FFE01D0007E01C00FAE01B000F";
attribute INIT_02 of ram_1024_x_18  : label is "E02A001FE0290000E028003FE0270000E026007FE0250000E02400FFE0230000";
attribute INIT_03 of ram_1024_x_18  : label is "E0320001E0310000E0300003E02F0000E02E0007E02D0000E02C000FE02B0000";
attribute INIT_04 of ram_1024_x_18  : label is "8001D01001130032EE090E01EE080E00ED390D00ED3A0D00EC370C74EC380C9B";
attribute INIT_05 of ram_1024_x_18  : label is "613750CDE90059A0EE08AEFF6E08EE098E006E09BEE00B130A100900E010000E";
attribute INIT_06 of ram_1024_x_18  : label is "020E507343001390623A6139E234E1335464C3010108020E5068430013906238";
attribute INIT_07 of ram_1024_x_18  : label is "03006409650806000700EF3B7F108101EF3C7F1011B0E236E135546FC3010108";
attribute INIT_08 of ram_1024_x_18  : label is "E03701660700060065366435030002006138603754A848010143000001000200";
attribute INIT_09 of ram_1024_x_18  : label is "0300020061086009E13AE039016B070006006534643303000200613A6039E138";
attribute INIT_0A of ram_1024_x_18  : label is "0700060065366435030002006138603740C9E108E009016607000600653C643B";
attribute INIT_0B of ram_1024_x_18  : label is "61086009E13AE0390166070006006534643303000200613A6039E138E037016B";
attribute INIT_0C of ram_1024_x_18  : label is "6038E00B6037405C8B018B018901E108E009016B07000600653C643B03000200";
attribute INIT_0D of ram_1024_x_18  : label is "0028010012600300013500D80109C201C302620B630AE00C603AE00D6039E00A";
attribute INIT_0E of ram_1024_x_18  : label is "603CE03B01700028010012600300013500220102C203C304620D630CE03C0170";
attribute INIT_0F of ram_1024_x_18  : label is "1170E000E10101221040116017301620151014004052C020003FC017603BC016";
attribute INIT_10 of ram_1024_x_18  : label is "66030700E006E107012210501170E004E105012210501160E002E10301221040";
attribute INIT_11 of ram_1024_x_18  : label is "0400050066066707016B6400650106000700016B000061046205030004006502";
attribute INIT_12 of ram_1024_x_18  : label is "113055280206040803089310512B3020040003000201E43DE33EE23FA000016B";
attribute INIT_13 of ram_1024_x_18  : label is "8601F510D40059425510E10054000600070014201530A000643D633E623F1040";
attribute INIT_14 of ram_1024_x_18  : label is "5400415B514F595955104163514B59615620415F5147595D5730A0004139A700";
attribute INIT_15 of ram_1024_x_18  : label is "0804416508014165080441650801416508044165080141650802415751535955";
attribute INIT_16 of ram_1024_x_18  : label is "A000B370B260B1509040A000F370F260F150D040A00041650804416508014165";
attribute INIT_17 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000004173A000B1309020";
attribute INIT_18 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_19 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "002182B6B40ADAD03992400A5088888888888888888888888888888888888888";
attribute INITP_01 of ram_1024_x_18 : label is "2B000E222C030A0B00C282222356B0000AC0002B0000EB0000AC0002B0000DC0";
attribute INITP_02 of ram_1024_x_18 : label is "000000E595655B333333333F7F7F7F6D575402003A9D02AB00C030000AC2B0AC";
attribute INITP_03 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A00D5E019001FE01800B6E017003EE01600B1E0150076E014000FE01300C9",
                INIT_01 => X"E02200FFE0210001E02000FFE01F0003E01E00FFE01D0007E01C00FAE01B000F",
                INIT_02 => X"E02A001FE0290000E028003FE0270000E026007FE0250000E02400FFE0230000",
                INIT_03 => X"E0320001E0310000E0300003E02F0000E02E0007E02D0000E02C000FE02B0000",
                INIT_04 => X"8001D01001130032EE090E01EE080E00ED390D00ED3A0D00EC370C74EC380C9B",
                INIT_05 => X"613750CDE90059A0EE08AEFF6E08EE098E006E09BEE00B130A100900E010000E",
                INIT_06 => X"020E507343001390623A6139E234E1335464C3010108020E5068430013906238",
                INIT_07 => X"03006409650806000700EF3B7F108101EF3C7F1011B0E236E135546FC3010108",
                INIT_08 => X"E03701660700060065366435030002006138603754A848010143000001000200",
                INIT_09 => X"0300020061086009E13AE039016B070006006534643303000200613A6039E138",
                INIT_0A => X"0700060065366435030002006138603740C9E108E009016607000600653C643B",
                INIT_0B => X"61086009E13AE0390166070006006534643303000200613A6039E138E037016B",
                INIT_0C => X"6038E00B6037405C8B018B018901E108E009016B07000600653C643B03000200",
                INIT_0D => X"0028010012600300013500D80109C201C302620B630AE00C603AE00D6039E00A",
                INIT_0E => X"603CE03B01700028010012600300013500220102C203C304620D630CE03C0170",
                INIT_0F => X"1170E000E10101221040116017301620151014004052C020003FC017603BC016",
                INIT_10 => X"66030700E006E107012210501170E004E105012210501160E002E10301221040",
                INIT_11 => X"0400050066066707016B6400650106000700016B000061046205030004006502",
                INIT_12 => X"113055280206040803089310512B3020040003000201E43DE33EE23FA000016B",
                INIT_13 => X"8601F510D40059425510E10054000600070014201530A000643D633E623F1040",
                INIT_14 => X"5400415B514F595955104163514B59615620415F5147595D5730A0004139A700",
                INIT_15 => X"0804416508014165080441650801416508044165080141650802415751535955",
                INIT_16 => X"A000B370B260B1509040A000F370F260F150D040A00041650804416508014165",
                INIT_17 => X"0000000000000000000000000000000000000000000000004173A000B1309020",
                INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"002182B6B40ADAD03992400A5088888888888888888888888888888888888888",
               INITP_01 => X"2B000E222C030A0B00C282222356B0000AC0002B0000EB0000AC0002B0000DC0",
               INITP_02 => X"000000E595655B333333333F7F7F7F6D575402003A9D02AB00C030000AC2B0AC",
               INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
