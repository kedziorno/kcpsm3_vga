--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A0003E01900FBE0180007E01700D7E016000EE01500D6E0140019E0130022";
attribute INIT_01 of ram_1024_x_18  : label is "E0220000E0210040E0200000E01F0080E01E0001E01D0000E01C0001E01B00FF";
attribute INIT_02 of ram_1024_x_18  : label is "E02A0000E0290004E0280000E0270008E0260000E0250010E0240000E0230020";
attribute INIT_03 of ram_1024_x_18  : label is "E00E0000E00D0000E00C0013E00B006FE02E0000E02D0001E02C0000E02B0002";
attribute INIT_04 of ram_1024_x_18  : label is "E031A0006031E03080016030E0310000E0300001E02F000E8001D0100113002E";
attribute INIT_05 of ram_1024_x_18  : label is "6001B0000500C003E0006031C003E0016030518A4404019F0068010162306331";
attribute INIT_06 of ram_1024_x_18  : label is "600F0503587DE010E0326010E00FE044600F05025886E010E032600FE001E044";
attribute INIT_07 of ram_1024_x_18  : label is "8001E0FF600FE010E0326010E00FE044600F05015886E010E0326010E00FE044";
attribute INIT_08 of ram_1024_x_18  : label is "E006000006000813E010A0326010E00F8044600F408CE010A000E0FF6010E00F";
attribute INIT_09 of ram_1024_x_18  : label is "04008801E01270808801E0117080E00A600EE009600DE008600CE007600B6706";
attribute INIT_0A of ram_1024_x_18  : label is "000A000A000AA08060101400D040000A000AA080600E1400D040000AA080600C";
attribute INIT_0B of ram_1024_x_18  : label is "6011E012A000E0FF6012E0118001E0FF601154BF4080A080601084011400D040";
attribute INIT_0C of ram_1024_x_18  : label is "0137012754D3C40140F40154013754CCC401E010B01061106012E00F9010610F";
attribute INIT_0D of ram_1024_x_18  : label is "C40140F4014B0137012F012754DFC40140F40137012F54D8C40140F40154014B";
attribute INIT_0E of ram_1024_x_18  : label is "40F40154014B0137012F54F0C40140F40137012754E9C40140F4014B013754E4";
attribute INIT_0F of ram_1024_x_18  : label is "E00D9010610D6007E00CB010610C600AE00B9010610B600901540137012F0127";
attribute INIT_10 of ram_1024_x_18  : label is "5126B05000034090410D550C56F06F2F8601E00680016006E00EB010610E6008";
attribute INIT_11 of ram_1024_x_18  : label is "E0FF600D5126B0500001E00CA000E0FF600CE00B8001E0FF600B511BB0500002";
attribute INIT_12 of ram_1024_x_18  : label is "B000A000E008E0006008E007E0016007B000415DE00EA000E0FF600EE00D8001";
attribute INIT_13 of ram_1024_x_18  : label is "6007E008000A6008B000C701514A50701070A000E00AE000600AE009E0016009";
attribute INIT_14 of ram_1024_x_18  : label is "6008E0078001E0FF6007A0004137E009000A6009E00A000A600AB000E007000A";
attribute INIT_15 of ram_1024_x_18  : label is "C002E003600BA000E00AA000E0FF600AE0098001E0FF6009A000E008A000E0FF";
attribute INIT_16 of ram_1024_x_18  : label is "019100330103C302C20262036302C001E004600EC001E005600DC002E002600C";
attribute INIT_17 of ram_1024_x_18  : label is "010012600300019100330103C301C20162056304E03C018E0028010012600300";
attribute INIT_18 of ram_1024_x_18  : label is "B1309020A000F130D020418A404AC020003FC017603BC016603CE03B018E0028";
attribute INIT_19 of ram_1024_x_18  : label is "5310A0004195A7008601F510D400599E5510E10054000600070014201530A000";
attribute INIT_1A of ram_1024_x_18  : label is "000000000000A000040441AC040241AC040141A955AB59A7520041AB51A359A7";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "42490E490E490E49028A370092488A5088888888888888888888888888888888";
attribute INITP_01 of ram_1024_x_18 : label is "909090FFFFF7FDFF7FFDFF7FFDFF642424243410A80280201862222080924E42";
attribute INITP_02 of ram_1024_x_18 : label is "030A0B00C2828A28A29090A4242E8A0A281D2924292439090C242430C3F46490";
attribute INITP_03 of ram_1024_x_18 : label is "000000000000000000000000000000000000000002333F7F6D575402597E222C";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A0003E01900FBE0180007E01700D7E016000EE01500D6E0140019E0130022",
                INIT_01 => X"E0220000E0210040E0200000E01F0080E01E0001E01D0000E01C0001E01B00FF",
                INIT_02 => X"E02A0000E0290004E0280000E0270008E0260000E0250010E0240000E0230020",
                INIT_03 => X"E00E0000E00D0000E00C0013E00B006FE02E0000E02D0001E02C0000E02B0002",
                INIT_04 => X"E031A0006031E03080016030E0310000E0300001E02F000E8001D0100113002E",
                INIT_05 => X"6001B0000500C003E0006031C003E0016030518A4404019F0068010162306331",
                INIT_06 => X"600F0503587DE010E0326010E00FE044600F05025886E010E032600FE001E044",
                INIT_07 => X"8001E0FF600FE010E0326010E00FE044600F05015886E010E0326010E00FE044",
                INIT_08 => X"E006000006000813E010A0326010E00F8044600F408CE010A000E0FF6010E00F",
                INIT_09 => X"04008801E01270808801E0117080E00A600EE009600DE008600CE007600B6706",
                INIT_0A => X"000A000A000AA08060101400D040000A000AA080600E1400D040000AA080600C",
                INIT_0B => X"6011E012A000E0FF6012E0118001E0FF601154BF4080A080601084011400D040",
                INIT_0C => X"0137012754D3C40140F40154013754CCC401E010B01061106012E00F9010610F",
                INIT_0D => X"C40140F4014B0137012F012754DFC40140F40137012F54D8C40140F40154014B",
                INIT_0E => X"40F40154014B0137012F54F0C40140F40137012754E9C40140F4014B013754E4",
                INIT_0F => X"E00D9010610D6007E00CB010610C600AE00B9010610B600901540137012F0127",
                INIT_10 => X"5126B05000034090410D550C56F06F2F8601E00680016006E00EB010610E6008",
                INIT_11 => X"E0FF600D5126B0500001E00CA000E0FF600CE00B8001E0FF600B511BB0500002",
                INIT_12 => X"B000A000E008E0006008E007E0016007B000415DE00EA000E0FF600EE00D8001",
                INIT_13 => X"6007E008000A6008B000C701514A50701070A000E00AE000600AE009E0016009",
                INIT_14 => X"6008E0078001E0FF6007A0004137E009000A6009E00A000A600AB000E007000A",
                INIT_15 => X"C002E003600BA000E00AA000E0FF600AE0098001E0FF6009A000E008A000E0FF",
                INIT_16 => X"019100330103C302C20262036302C001E004600EC001E005600DC002E002600C",
                INIT_17 => X"010012600300019100330103C301C20162056304E03C018E0028010012600300",
                INIT_18 => X"B1309020A000F130D020418A404AC020003FC017603BC016603CE03B018E0028",
                INIT_19 => X"5310A0004195A7008601F510D400599E5510E10054000600070014201530A000",
                INIT_1A => X"000000000000A000040441AC040241AC040141A955AB59A7520041AB51A359A7",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"42490E490E490E49028A370092488A5088888888888888888888888888888888",
               INITP_01 => X"909090FFFFF7FDFF7FFDFF7FFDFF642424243410A80280201862222080924E42",
               INITP_02 => X"030A0B00C2828A28A29090A4242E8A0A281D2924292439090C242430C3F46490",
               INITP_03 => X"000000000000000000000000000000000000000002333F7F6D575402597E222C",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
