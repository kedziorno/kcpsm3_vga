--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A0003E01900FBE0180007E01700D7E016000EE01500D6E0140019E0130022";
attribute INIT_01 of ram_1024_x_18  : label is "E0220000E0210040E0200000E01F0080E01E0001E01D0000E01C0001E01B00FF";
attribute INIT_02 of ram_1024_x_18  : label is "E02A0000E0290004E0280000E0270008E0260000E0250010E0240000E0230020";
attribute INIT_03 of ram_1024_x_18  : label is "E00E0000E00D0000E00C0013E00B006FE02E0000E02D0001E02C0000E02B0002";
attribute INIT_04 of ram_1024_x_18  : label is "0060E031008CE0300009E0310000E0300000E02F000E8001D0100113002E0500";
attribute INIT_05 of ram_1024_x_18  : label is "41A70060E03100C9E03000100060E0310010E03000C90060E0310009E030008C";
attribute INIT_06 of ram_1024_x_18  : label is "0502588FE010E032600FE001E0446001B0000500C003E0006031C003E0016030";
attribute INIT_07 of ram_1024_x_18  : label is "0501588FE010E0326010E00FE044600F05035886E010E0326010E00FE044600F";
attribute INIT_08 of ram_1024_x_18  : label is "600F4095E010A000E0FF6010E00F8001E0FF600FE010E0326010E00FE044600F";
attribute INIT_09 of ram_1024_x_18  : label is "E009600DE008600CE007600B6706E006000006000813E010A0326010E00F8044";
attribute INIT_0A of ram_1024_x_18  : label is "A080600E1400D0400000A080600C04008801E01270808801E0117080E00A600E";
attribute INIT_0B of ram_1024_x_18  : label is "4000B0106110008084011400D040000000000000A08060101400D04000000000";
attribute INIT_0C of ram_1024_x_18  : label is "B01061106012E00F9010610F6011E012A000E0FF6012E0118001E0FF601154C9";
attribute INIT_0D of ram_1024_x_18  : label is "C40141050168015F014B013B54DF4400C40141050168014B54D74400C401E010";
attribute INIT_0E of ram_1024_x_18  : label is "54F34400C4014105015F014B0143013B54ED4400C4014105014B014354E54400";
attribute INIT_0F of ram_1024_x_18  : label is "0168015F014B014355014400C4014105014B013B54F94400C4014105015F014B";
attribute INIT_10 of ram_1024_x_18  : label is "9010610D6007E00CB010610C600AE00B9010610B60090168014B0143013B4105";
attribute INIT_11 of ram_1024_x_18  : label is "B05000034099411E551D56F06F2F8601E00680016006E00EB010610E6008E00D";
attribute INIT_12 of ram_1024_x_18  : label is "B0500001E00CA000E0FF600CE00B8001E0FF600B512E4000B0500002513A4000";
attribute INIT_13 of ram_1024_x_18  : label is "6008E007E0016007B0004171E00EA000E0FF600EE00D8001E0FF600D513A4000";
attribute INIT_14 of ram_1024_x_18  : label is "B000C701515E40001070A000E00AE000600AE009E0016009B000A000E008E000";
attribute INIT_15 of ram_1024_x_18  : label is "6007A000414BE009000A6009E00A000A600AB000E007000A6007E008000A6008";
attribute INIT_16 of ram_1024_x_18  : label is "E00AA000E0FF600AE0098001E0FF6009A000E008A000E0FF6008E0078001E0FF";
attribute INIT_17 of ram_1024_x_18  : label is "6003C0026002C0026002C0026003E004600EE005600DE002600CE003600BA000";
attribute INIT_18 of ram_1024_x_18  : label is "030001AE0033010362026303A000C0016005C0016004C0016004C0016005C002";
attribute INIT_19 of ram_1024_x_18  : label is "E03B01AB002801001260030001AE0033010362046305E03C01AB002801001260";
attribute INIT_1A of ram_1024_x_18  : label is "14201530A000B1309020A000F130D02041A7404BC020003FC017603BC016603C";
attribute INIT_1B of ram_1024_x_18  : label is "41C851C059C45310A00041B2A7008601F510D40059BB5510E100540006000700";
attribute INIT_1C of ram_1024_x_18  : label is "000000000000000000000000A000040441C9040241C9040141C655C859C45200";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "3924392439240A28F88E2388E222294088888888888888888888888888888888";
attribute INITP_01 of ram_1024_x_18 : label is "FFD7FD7FD7FFD7FD7FFD7FD6424242434042A00A008061888882024939090924";
attribute INITP_02 of ram_1024_x_18 : label is "222222229090A4242E8A0A281D2924292439090D09090D0D0FD19242424243FF";
attribute INITP_03 of ram_1024_x_18 : label is "0000000000000000000000000008CCFDFDB55D500965F888B00C02C0300A2222";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A0003E01900FBE0180007E01700D7E016000EE01500D6E0140019E0130022",
                INIT_01 => X"E0220000E0210040E0200000E01F0080E01E0001E01D0000E01C0001E01B00FF",
                INIT_02 => X"E02A0000E0290004E0280000E0270008E0260000E0250010E0240000E0230020",
                INIT_03 => X"E00E0000E00D0000E00C0013E00B006FE02E0000E02D0001E02C0000E02B0002",
                INIT_04 => X"0060E031008CE0300009E0310000E0300000E02F000E8001D0100113002E0500",
                INIT_05 => X"41A70060E03100C9E03000100060E0310010E03000C90060E0310009E030008C",
                INIT_06 => X"0502588FE010E032600FE001E0446001B0000500C003E0006031C003E0016030",
                INIT_07 => X"0501588FE010E0326010E00FE044600F05035886E010E0326010E00FE044600F",
                INIT_08 => X"600F4095E010A000E0FF6010E00F8001E0FF600FE010E0326010E00FE044600F",
                INIT_09 => X"E009600DE008600CE007600B6706E006000006000813E010A0326010E00F8044",
                INIT_0A => X"A080600E1400D0400000A080600C04008801E01270808801E0117080E00A600E",
                INIT_0B => X"4000B0106110008084011400D040000000000000A08060101400D04000000000",
                INIT_0C => X"B01061106012E00F9010610F6011E012A000E0FF6012E0118001E0FF601154C9",
                INIT_0D => X"C40141050168015F014B013B54DF4400C40141050168014B54D74400C401E010",
                INIT_0E => X"54F34400C4014105015F014B0143013B54ED4400C4014105014B014354E54400",
                INIT_0F => X"0168015F014B014355014400C4014105014B013B54F94400C4014105015F014B",
                INIT_10 => X"9010610D6007E00CB010610C600AE00B9010610B60090168014B0143013B4105",
                INIT_11 => X"B05000034099411E551D56F06F2F8601E00680016006E00EB010610E6008E00D",
                INIT_12 => X"B0500001E00CA000E0FF600CE00B8001E0FF600B512E4000B0500002513A4000",
                INIT_13 => X"6008E007E0016007B0004171E00EA000E0FF600EE00D8001E0FF600D513A4000",
                INIT_14 => X"B000C701515E40001070A000E00AE000600AE009E0016009B000A000E008E000",
                INIT_15 => X"6007A000414BE009000A6009E00A000A600AB000E007000A6007E008000A6008",
                INIT_16 => X"E00AA000E0FF600AE0098001E0FF6009A000E008A000E0FF6008E0078001E0FF",
                INIT_17 => X"6003C0026002C0026002C0026003E004600EE005600DE002600CE003600BA000",
                INIT_18 => X"030001AE0033010362026303A000C0016005C0016004C0016004C0016005C002",
                INIT_19 => X"E03B01AB002801001260030001AE0033010362046305E03C01AB002801001260",
                INIT_1A => X"14201530A000B1309020A000F130D02041A7404BC020003FC017603BC016603C",
                INIT_1B => X"41C851C059C45310A00041B2A7008601F510D40059BB5510E100540006000700",
                INIT_1C => X"000000000000000000000000A000040441C9040241C9040141C655C859C45200",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"3924392439240A28F88E2388E222294088888888888888888888888888888888",
               INITP_01 => X"FFD7FD7FD7FFD7FD7FFD7FD6424242434042A00A008061888882024939090924",
               INITP_02 => X"222222229090A4242E8A0A281D2924292439090D09090D0D0FD19242424243FF",
               INITP_03 => X"0000000000000000000000000008CCFDFDB55D500965F888B00C02C0300A2222",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
