--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A00D5E019001FE01800B6E017003EE01600B1E0150076E014000FE01300C9";
attribute INIT_01 of ram_1024_x_18  : label is "E02200FFE0210001E02000FFE01F0003E01E00FFE01D0007E01C00FAE01B000F";
attribute INIT_02 of ram_1024_x_18  : label is "E02A001FE0290000E028003FE0270000E026007FE0250000E02400FFE0230000";
attribute INIT_03 of ram_1024_x_18  : label is "E0320001E0310000E0300003E02F0000E02E0007E02D0000E02C000FE02B0000";
attribute INIT_04 of ram_1024_x_18  : label is "8001D01001130032EE3D0E01EE3E0E00ED390D00ED3A0D00EC370C9BEC380C74";
attribute INIT_05 of ram_1024_x_18  : label is "50CF59A0EE3EAE04CE036E3EEE3D8E77CE036E3DBEE00B130A0F0900E010000E";
attribute INIT_06 of ram_1024_x_18  : label is "507443001390623A6139E234E1335465C3010108020E50694300139062386137";
attribute INIT_07 of ram_1024_x_18  : label is "EF086F3EEF096F3DEF3B7F108101EF3C7F1011B0E236E1355470C3010108020E";
attribute INIT_08 of ram_1024_x_18  : label is "0700060065366435030002006138603754AAA380A300E3FF63088201E2FF6209";
attribute INIT_09 of ram_1024_x_18  : label is "61086009E13AE039016D070006006534643303000200613A6039E138E0370168";
attribute INIT_0A of ram_1024_x_18  : label is "65366435030002006138603740CBE108E009016807000600653C643B03000200";
attribute INIT_0B of ram_1024_x_18  : label is "E13AE0390168070006006534643303000200613A6039E138E037016D07000600";
attribute INIT_0C of ram_1024_x_18  : label is "6037405E8B018B018901E108E009016D07000600653C643B0300020061086009";
attribute INIT_0D of ram_1024_x_18  : label is "12600300013700D80109C302C202620B630AE00C603AE00D6039E00A6038E00B";
attribute INIT_0E of ram_1024_x_18  : label is "0172002801A912600300013700220102C301C201620D630CE03C017200280100";
attribute INIT_0F of ram_1024_x_18  : label is "E10101241040116017301620151014004052C020003FC017603BC016603CE03B";
attribute INIT_10 of ram_1024_x_18  : label is "E006E107012410501170E004E105012410501160E002E103012410401170E000";
attribute INIT_11 of ram_1024_x_18  : label is "66066707016D6400650106000700016D00006104620503000400650266030700";
attribute INIT_12 of ram_1024_x_18  : label is "0206040803089310512D3020040003000201E43DE33EE23FA000016D04000500";
attribute INIT_13 of ram_1024_x_18  : label is "D40059445510E10054000600070014201530A000643D633E623F10401130552A";
attribute INIT_14 of ram_1024_x_18  : label is "5151595B55104165514D5963562041615149595F5730A000413BA7008601F510";
attribute INIT_15 of ram_1024_x_18  : label is "080141670804416708014167080441670801416708024159515559575400415D";
attribute INIT_16 of ram_1024_x_18  : label is "B260B1509040A000F370F260F150D040A0004167080441670801416708044167";
attribute INIT_17 of ram_1024_x_18  : label is "040241820401417F5581597D520041815179597D5310A000B1309020A000B370";
attribute INIT_18 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000004183A00004044182";
attribute INIT_19 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "88860ADAD02B6B40D989800A5088888888888888888888888888888888888888";
attribute INITP_01 of ram_1024_x_18 : label is "B000E222C030A0B00C282222356B0000AC0002B0000EB0000AC0002B0000C410";
attribute INITP_02 of ram_1024_x_18 : label is "33F7F6595655B333333333F7F7F7F6D575402003A9D02AB00C030000AC2B0AC2";
attribute INITP_03 of ram_1024_x_18 : label is "00000000000000000000000000000000000000000000000000000000000000E3";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A00D5E019001FE01800B6E017003EE01600B1E0150076E014000FE01300C9",
                INIT_01 => X"E02200FFE0210001E02000FFE01F0003E01E00FFE01D0007E01C00FAE01B000F",
                INIT_02 => X"E02A001FE0290000E028003FE0270000E026007FE0250000E02400FFE0230000",
                INIT_03 => X"E0320001E0310000E0300003E02F0000E02E0007E02D0000E02C000FE02B0000",
                INIT_04 => X"8001D01001130032EE3D0E01EE3E0E00ED390D00ED3A0D00EC370C9BEC380C74",
                INIT_05 => X"50CF59A0EE3EAE04CE036E3EEE3D8E77CE036E3DBEE00B130A0F0900E010000E",
                INIT_06 => X"507443001390623A6139E234E1335465C3010108020E50694300139062386137",
                INIT_07 => X"EF086F3EEF096F3DEF3B7F108101EF3C7F1011B0E236E1355470C3010108020E",
                INIT_08 => X"0700060065366435030002006138603754AAA380A300E3FF63088201E2FF6209",
                INIT_09 => X"61086009E13AE039016D070006006534643303000200613A6039E138E0370168",
                INIT_0A => X"65366435030002006138603740CBE108E009016807000600653C643B03000200",
                INIT_0B => X"E13AE0390168070006006534643303000200613A6039E138E037016D07000600",
                INIT_0C => X"6037405E8B018B018901E108E009016D07000600653C643B0300020061086009",
                INIT_0D => X"12600300013700D80109C302C202620B630AE00C603AE00D6039E00A6038E00B",
                INIT_0E => X"0172002801A912600300013700220102C301C201620D630CE03C017200280100",
                INIT_0F => X"E10101241040116017301620151014004052C020003FC017603BC016603CE03B",
                INIT_10 => X"E006E107012410501170E004E105012410501160E002E103012410401170E000",
                INIT_11 => X"66066707016D6400650106000700016D00006104620503000400650266030700",
                INIT_12 => X"0206040803089310512D3020040003000201E43DE33EE23FA000016D04000500",
                INIT_13 => X"D40059445510E10054000600070014201530A000643D633E623F10401130552A",
                INIT_14 => X"5151595B55104165514D5963562041615149595F5730A000413BA7008601F510",
                INIT_15 => X"080141670804416708014167080441670801416708024159515559575400415D",
                INIT_16 => X"B260B1509040A000F370F260F150D040A0004167080441670801416708044167",
                INIT_17 => X"040241820401417F5581597D520041815179597D5310A000B1309020A000B370",
                INIT_18 => X"0000000000000000000000000000000000000000000000004183A00004044182",
                INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"88860ADAD02B6B40D989800A5088888888888888888888888888888888888888",
               INITP_01 => X"B000E222C030A0B00C282222356B0000AC0002B0000EB0000AC0002B0000C410",
               INITP_02 => X"33F7F6595655B333333333F7F7F7F6D575402003A9D02AB00C030000AC2B0AC2",
               INITP_03 => X"00000000000000000000000000000000000000000000000000000000000000E3",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
