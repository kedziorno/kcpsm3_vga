--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E91A0903E91909FBE9180907E91709D7E916090EE91509D6E9140919E9130922";
attribute INIT_01 of ram_1024_x_18  : label is "E9220900E9210940E9200900E91F0980E91E0901E91D0900E91C0901E91B09FF";
attribute INIT_02 of ram_1024_x_18  : label is "E92A0900E9290904E9280900E9270908E9260900E9250910E9240900E9230920";
attribute INIT_03 of ram_1024_x_18  : label is "E90E0900E90D0900E90C0913E90B096FE92E0900E92D0901E92C0900E92B0902";
attribute INIT_04 of ram_1024_x_18  : label is "C9170977C916099FC920093FC9170900C9160900E92F090E8901D9100113092E";
attribute INIT_05 of ram_1024_x_18  : label is "0FD70EB2C920093FC9170977C9160900C920093FC9170900C916099FC920093F";
attribute INIT_06 of ram_1024_x_18  : label is "C201C302620363020095EF00EE0151FE4404019E10E011F0024E0328AF008E39";
attribute INIT_07 of ram_1024_x_18  : label is "C30462056304E03C01EB0028010002000300060007001460157001F000330103";
attribute INIT_08 of ram_1024_x_18  : label is "C916693CE03B01EB0028010002000300060007001460157001F000330103C203";
attribute INIT_09 of ram_1024_x_18  : label is "690F060258BEE910E9326900E90FE9446901B99006004060C920093FC917693B";
attribute INIT_0A of ram_1024_x_18  : label is "690F060158BEE910E9326910E90FE944690F060358B5E910E9326910E90FE944";
attribute INIT_0B of ram_1024_x_18  : label is "8944690F40C4E910A900E9FF6910E90F8901E9FF690FE910E9326910E90FE944";
attribute INIT_0C of ram_1024_x_18  : label is "690EE909690DE908690CE907690B6406E906090005000A13E910A9326910E90F";
attribute INIT_0D of ram_1024_x_18  : label is "690E1790D970090EA980690C07008A018A01E91279B08B01E91179B01BA0E90A";
attribute INIT_0E of ram_1024_x_18  : label is "54F8A980691087011790D970090E090E090EA98069101790D970090E090EA980";
attribute INIT_0F of ram_1024_x_18  : label is "E910B91061106912E90F9910610F6911E912A900E9FF6912E9118901E9FF6911";
attribute INIT_10 of ram_1024_x_18  : label is "017001685511C701412D018C018301700160550CC701412D018C01705505C701";
attribute INIT_11 of ram_1024_x_18  : label is "01605522C701412D01830170551DC701412D01830170016801605518C701412D";
attribute INIT_12 of ram_1024_x_18  : label is "9910610B6909018C017001680160412D018C0183017001685529C701412D0170";
attribute INIT_13 of ram_1024_x_18  : label is "E90689016906E90EB910610E6908E90D9910610D6907E90CB910610C690AE90B";
attribute INIT_14 of ram_1024_x_18  : label is "E90B8901E9FF690B5154B9600902515FB960090340C8414655455590692F8501";
attribute INIT_15 of ram_1024_x_18  : label is "4195E90EA900E9FF690EE90D8901E9FF690D515FB9600901E90CA900E9FF690C";
attribute INIT_16 of ram_1024_x_18  : label is "A000E90AE900690AE909E9016909B990A000E908E9006908E907E9016907B990";
attribute INIT_17 of ram_1024_x_18  : label is "09086909E90A0908690AB990E90709086907E90809086908B990C40151821940";
attribute INIT_18 of ram_1024_x_18  : label is "E9098901E9FF6909A000E908A900E9FF6908E9078901E9FF6907A0004170E909";
attribute INIT_19 of ram_1024_x_18  : label is "59A65310A000E904690EE905690DE902690CE903690BA000E90AA900E9FF690A";
attribute INIT_1A of ram_1024_x_18  : label is "1730162015101400A000040441AB040241AB040141A855AA59A6520041AA51A2";
attribute INIT_1B of ram_1024_x_18  : label is "1170E004E10501D810501160E002E10301D810401170E000E10101D810401160";
attribute INIT_1C of ram_1024_x_18  : label is "65010600070001EB00006104620503000400650266030700E006E10701D81050";
attribute INIT_1D of ram_1024_x_18  : label is "51E13020040003000201E43DE33EE23FA00001EB040005006606670701EB6400";
attribute INIT_1E of ram_1024_x_18  : label is "A000B370B260B1509040A000643D633E623F1040113055DE0206040803089310";
attribute INIT_1F of ram_1024_x_18  : label is "41FF41FFA00041F4A7008601F510D40059FD5510E10054000600070014201530";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "82C00030A0EB70050888888888888A5088888888888888888888888888888888";
attribute INITP_01 of ram_1024_x_18 : label is "90909090C10A802802016182222080924E4242490E490E490E4903888B0000C2";
attribute INITP_02 of ram_1024_x_18 : label is "8A0A281CA490A490E424309090C30FD19242424243FFFFDFF7FDFFF7FDFFF7FD";
attribute INITP_03 of ram_1024_x_18 : label is "FB55D500956003A9D02AB00C030000AC2B0AC2B0008CCFDFDA22229090A4242E";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E91A0903E91909FBE9180907E91709D7E916090EE91509D6E9140919E9130922",
                INIT_01 => X"E9220900E9210940E9200900E91F0980E91E0901E91D0900E91C0901E91B09FF",
                INIT_02 => X"E92A0900E9290904E9280900E9270908E9260900E9250910E9240900E9230920",
                INIT_03 => X"E90E0900E90D0900E90C0913E90B096FE92E0900E92D0901E92C0900E92B0902",
                INIT_04 => X"C9170977C916099FC920093FC9170900C9160900E92F090E8901D9100113092E",
                INIT_05 => X"0FD70EB2C920093FC9170977C9160900C920093FC9170900C916099FC920093F",
                INIT_06 => X"C201C302620363020095EF00EE0151FE4404019E10E011F0024E0328AF008E39",
                INIT_07 => X"C30462056304E03C01EB0028010002000300060007001460157001F000330103",
                INIT_08 => X"C916693CE03B01EB0028010002000300060007001460157001F000330103C203",
                INIT_09 => X"690F060258BEE910E9326900E90FE9446901B99006004060C920093FC917693B",
                INIT_0A => X"690F060158BEE910E9326910E90FE944690F060358B5E910E9326910E90FE944",
                INIT_0B => X"8944690F40C4E910A900E9FF6910E90F8901E9FF690FE910E9326910E90FE944",
                INIT_0C => X"690EE909690DE908690CE907690B6406E906090005000A13E910A9326910E90F",
                INIT_0D => X"690E1790D970090EA980690C07008A018A01E91279B08B01E91179B01BA0E90A",
                INIT_0E => X"54F8A980691087011790D970090E090E090EA98069101790D970090E090EA980",
                INIT_0F => X"E910B91061106912E90F9910610F6911E912A900E9FF6912E9118901E9FF6911",
                INIT_10 => X"017001685511C701412D018C018301700160550CC701412D018C01705505C701",
                INIT_11 => X"01605522C701412D01830170551DC701412D01830170016801605518C701412D",
                INIT_12 => X"9910610B6909018C017001680160412D018C0183017001685529C701412D0170",
                INIT_13 => X"E90689016906E90EB910610E6908E90D9910610D6907E90CB910610C690AE90B",
                INIT_14 => X"E90B8901E9FF690B5154B9600902515FB960090340C8414655455590692F8501",
                INIT_15 => X"4195E90EA900E9FF690EE90D8901E9FF690D515FB9600901E90CA900E9FF690C",
                INIT_16 => X"A000E90AE900690AE909E9016909B990A000E908E9006908E907E9016907B990",
                INIT_17 => X"09086909E90A0908690AB990E90709086907E90809086908B990C40151821940",
                INIT_18 => X"E9098901E9FF6909A000E908A900E9FF6908E9078901E9FF6907A0004170E909",
                INIT_19 => X"59A65310A000E904690EE905690DE902690CE903690BA000E90AA900E9FF690A",
                INIT_1A => X"1730162015101400A000040441AB040241AB040141A855AA59A6520041AA51A2",
                INIT_1B => X"1170E004E10501D810501160E002E10301D810401170E000E10101D810401160",
                INIT_1C => X"65010600070001EB00006104620503000400650266030700E006E10701D81050",
                INIT_1D => X"51E13020040003000201E43DE33EE23FA00001EB040005006606670701EB6400",
                INIT_1E => X"A000B370B260B1509040A000643D633E623F1040113055DE0206040803089310",
                INIT_1F => X"41FF41FFA00041F4A7008601F510D40059FD5510E10054000600070014201530",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"82C00030A0EB70050888888888888A5088888888888888888888888888888888",
               INITP_01 => X"90909090C10A802802016182222080924E4242490E490E490E4903888B0000C2",
               INITP_02 => X"8A0A281CA490A490E424309090C30FD19242424243FFFFDFF7FDFFF7FDFFF7FD",
               INITP_03 => X"FB55D500956003A9D02AB00C030000AC2B0AC2B0008CCFDFDA22229090A4242E",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
