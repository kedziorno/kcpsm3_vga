--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A0000E0190001E0180001E0170003E0160005E015000AE0140013E0130020";
attribute INIT_01 of ram_1024_x_18  : label is "0A080900ED390D00EC370C4DE010000E8001D0100113001AEE3D0E00EE3E0E00";
attribute INIT_02 of ram_1024_x_18  : label is "515A4201623E4062502D4268623DEE3EAE00CE036E3EEE3D8E01CE036E3D0B13";
attribute INIT_03 of ram_1024_x_18  : label is "0300E024000254474401014C00B40100623D633E4062E02400015436405A603D";
attribute INIT_04 of ram_1024_x_18  : label is "E024000354584401014C000E0101623D633E4062E03DE13E010B603D613E02B4";
attribute INIT_05 of ram_1024_x_18  : label is "E2FF623EE23D8201E2FF623DE02400044062E03DE13E010B00B40100023D033E";
attribute INIT_06 of ram_1024_x_18  : label is "E133546CC301010A506F43001390613750A159A0EF086F3EEF096F3DE23EA200";
attribute INIT_07 of ram_1024_x_18  : label is "6037508F4480A4806408EF3B7F1011B0E1355474C301010A5077430013906139";
attribute INIT_08 of ram_1024_x_18  : label is "6037409EE108E009E100D020623B61086009E039904064336039E037D0406435";
attribute INIT_09 of ram_1024_x_18  : label is "8B018901E108E009A1009020623B61086009E039D04064336039E03790406435";
attribute INIT_0A of ram_1024_x_18  : label is "400250B24001602440B7E0378001E0FF603740AC50A7400450A7400160244066";
attribute INIT_0B of ram_1024_x_18  : label is "E0228028000AC001600DE00D6039E00B603740B7E0398001E0FF603940B750B2";
attribute INIT_0C of ram_1024_x_18  : label is "1730162015101400401AC020003FC0176023C0166022E0238028000AC002600B";
attribute INIT_0D of ram_1024_x_18  : label is "1170E004E10500F810501160E002E10300F810401170E000E10100F810401160";
attribute INIT_0E of ram_1024_x_18  : label is "650106000700014400006104620503000400650266030700E006E10700F81050";
attribute INIT_0F of ram_1024_x_18  : label is "51013020040003000201E43DE33EE23FA0000144040005006606670701446400";
attribute INIT_10 of ram_1024_x_18  : label is "14201530A000F130D020A000643D633E623F1040113054FE0206040803089310";
attribute INIT_11 of ram_1024_x_18  : label is "4138512059365730A0004112A7008601F510D400591B5510E100540006000700";
attribute INIT_12 of ram_1024_x_18  : label is "413E0801413E08024130512C592E54004134512859325510413C5124593A5620";
attribute INIT_13 of ram_1024_x_18  : label is "D040A000413E0804413E0801413E0804413E0801413E0804413E0801413E0804";
attribute INIT_14 of ram_1024_x_18  : label is "4158515059545310A000B1309020A000B370B260B1509040A000F370F260F150";
attribute INIT_15 of ram_1024_x_18  : label is "00000000000000000000415AA000040441590402415904014156555859545200";
attribute INIT_16 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_17 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_18 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_19 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "3420B6D0B6D0D8890908EB008DC03AC023700E34D3D26260088A508888888888";
attribute INITP_01 of ram_1024_x_18 : label is "D02AB00C030000AC2B0AC2B000E222689A22390F74E43DD35A5024243A502424";
attribute INITP_02 of ram_1024_x_18 : label is "00000000000000000038CCFDFD9655956CCCCCCCCCFDFDFDFDB55D50096003A9";
attribute INITP_03 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A0000E0190001E0180001E0170003E0160005E015000AE0140013E0130020",
                INIT_01 => X"0A080900ED390D00EC370C4DE010000E8001D0100113001AEE3D0E00EE3E0E00",
                INIT_02 => X"515A4201623E4062502D4268623DEE3EAE00CE036E3EEE3D8E01CE036E3D0B13",
                INIT_03 => X"0300E024000254474401014C00B40100623D633E4062E02400015436405A603D",
                INIT_04 => X"E024000354584401014C000E0101623D633E4062E03DE13E010B603D613E02B4",
                INIT_05 => X"E2FF623EE23D8201E2FF623DE02400044062E03DE13E010B00B40100023D033E",
                INIT_06 => X"E133546CC301010A506F43001390613750A159A0EF086F3EEF096F3DE23EA200",
                INIT_07 => X"6037508F4480A4806408EF3B7F1011B0E1355474C301010A5077430013906139",
                INIT_08 => X"6037409EE108E009E100D020623B61086009E039904064336039E037D0406435",
                INIT_09 => X"8B018901E108E009A1009020623B61086009E039D04064336039E03790406435",
                INIT_0A => X"400250B24001602440B7E0378001E0FF603740AC50A7400450A7400160244066",
                INIT_0B => X"E0228028000AC001600DE00D6039E00B603740B7E0398001E0FF603940B750B2",
                INIT_0C => X"1730162015101400401AC020003FC0176023C0166022E0238028000AC002600B",
                INIT_0D => X"1170E004E10500F810501160E002E10300F810401170E000E10100F810401160",
                INIT_0E => X"650106000700014400006104620503000400650266030700E006E10700F81050",
                INIT_0F => X"51013020040003000201E43DE33EE23FA0000144040005006606670701446400",
                INIT_10 => X"14201530A000F130D020A000643D633E623F1040113054FE0206040803089310",
                INIT_11 => X"4138512059365730A0004112A7008601F510D400591B5510E100540006000700",
                INIT_12 => X"413E0801413E08024130512C592E54004134512859325510413C5124593A5620",
                INIT_13 => X"D040A000413E0804413E0801413E0804413E0801413E0804413E0801413E0804",
                INIT_14 => X"4158515059545310A000B1309020A000B370B260B1509040A000F370F260F150",
                INIT_15 => X"00000000000000000000415AA000040441590402415904014156555859545200",
                INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"3420B6D0B6D0D8890908EB008DC03AC023700E34D3D26260088A508888888888",
               INITP_01 => X"D02AB00C030000AC2B0AC2B000E222689A22390F74E43DD35A5024243A502424",
               INITP_02 => X"00000000000000000038CCFDFD9655956CCCCCCCCCFDFDFDFDB55D50096003A9",
               INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
