--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A0003E01900FBE0180007E01700D7E016000EE01500D6E0140019E0130022";
attribute INIT_01 of ram_1024_x_18  : label is "E0220000E0210040E0200000E01F0080E01E0001E01D0000E01C0001E01B00FF";
attribute INIT_02 of ram_1024_x_18  : label is "E02A0000E0290004E0280000E0270008E0260000E0250010E0240000E0230020";
attribute INIT_03 of ram_1024_x_18  : label is "E00E0000E00D0000E00C0013E00B006FE02E0000E02D0001E02C0000E02B0002";
attribute INIT_04 of ram_1024_x_18  : label is "0060E031008CE0300009E0310000E0300000E02F000E8001D0100113002E0500";
attribute INIT_05 of ram_1024_x_18  : label is "41B30060E03100C9E03000100060E0310010E03000C90060E0310009E030008C";
attribute INIT_06 of ram_1024_x_18  : label is "0502588FE110E00FE132C04461006001B0000500C005E0006031C005E0016030";
attribute INIT_07 of ram_1024_x_18  : label is "0501588FE110E00FE132C0446110600F05035886E110E00FE132C0446110600F";
attribute INIT_08 of ram_1024_x_18  : label is "600F4095E010A000E0FF6010E00F8001E0FF600FE110E00FE132C0446110600F";
attribute INIT_09 of ram_1024_x_18  : label is "E009600DE008600CE007600B6706E006000006000813E110E00FA13280446110";
attribute INIT_0A of ram_1024_x_18  : label is "0002A080600C0400C207C106621261118801E01270808801E0117080E00A600E";
attribute INIT_0B of ram_1024_x_18  : label is "84011400D040000200020002A08060101400D04000020002A080600E1400D040";
attribute INIT_0C of ram_1024_x_18  : label is "C10662126111E012A000E0FF6012E0118001E0FF601150D12080B01001806010";
attribute INIT_0D of ram_1024_x_18  : label is "54E34400C401C0050010C005000FE010B01061106012E00F9010610F6011C207";
attribute INIT_0E of ram_1024_x_18  : label is "0157014F54F14400C40141110174016B0157014754EB4400C401411101740157";
attribute INIT_0F of ram_1024_x_18  : label is "C4014111016B015754FF4400C4014111016B0157014F014754F94400C4014111";
attribute INIT_10 of ram_1024_x_18  : label is "0157014F014741110174016B0157014F550D4400C40141110157014755054400";
attribute INIT_11 of ram_1024_x_18  : label is "E00DB130902063086207610E600DE10CE00BB1309020630A6209610C600B0174";
attribute INIT_12 of ram_1024_x_18  : label is "B050000251464000B05000034099412A552956F06F2F8601E00680016006E10E";
attribute INIT_13 of ram_1024_x_18  : label is "E0FF600D51464000B0500001E00CA000E0FF600CE00B8001E0FF600B513A4000";
attribute INIT_14 of ram_1024_x_18  : label is "B000A000E008E0006008E007E0016007B000417DE00EA000E0FF600EE00D8001";
attribute INIT_15 of ram_1024_x_18  : label is "6007E008000A6008B000C701516A40001070A000E00AE000600AE009E0016009";
attribute INIT_16 of ram_1024_x_18  : label is "6008E0078001E0FF6007A0004157E00900086009E00A000A600AB000E0070008";
attribute INIT_17 of ram_1024_x_18  : label is "600CE003600BA000E00AA000E0FF600AE0098001E0FF6009A000E008A000E0FF";
attribute INIT_18 of ram_1024_x_18  : label is "6004C0016005C0046003C0046002C0026002C0026003E004600EE005600DE002";
attribute INIT_19 of ram_1024_x_18  : label is "01B7002801001260030001BA0033010362026303A000C0036005C0036004C001";
attribute INIT_1A of ram_1024_x_18  : label is "C017603BC016603CE03B01B7002801001260030001BA0033010362046305E03C";
attribute INIT_1B of ram_1024_x_18  : label is "E10054000600070014201530A000B1309020A000F130D02041B3404BC020003F";
attribute INIT_1C of ram_1024_x_18  : label is "41D255D459D0520041D451CC59D05310A00041BEA7008601F510D40059C75510";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000A000040441D5040241D50401";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "3A503A503A500A28F88E2388E222294088888888888888888888888888888888";
attribute INITP_01 of ram_1024_x_18 : label is "7FD7FFD7FD7FFD7FD62242428242434042A00A0080A061888882029439090A50";
attribute INITP_02 of ram_1024_x_18 : label is "229090A4242E8A0A281D2924292439090D09090D0D0FD19294029403FFFFD7FD";
attribute INITP_03 of ram_1024_x_18 : label is "0000000000000000000008CCFDFDB55D500965F888B00C02C0300A2222222222";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A0003E01900FBE0180007E01700D7E016000EE01500D6E0140019E0130022",
                INIT_01 => X"E0220000E0210040E0200000E01F0080E01E0001E01D0000E01C0001E01B00FF",
                INIT_02 => X"E02A0000E0290004E0280000E0270008E0260000E0250010E0240000E0230020",
                INIT_03 => X"E00E0000E00D0000E00C0013E00B006FE02E0000E02D0001E02C0000E02B0002",
                INIT_04 => X"0060E031008CE0300009E0310000E0300000E02F000E8001D0100113002E0500",
                INIT_05 => X"41B30060E03100C9E03000100060E0310010E03000C90060E0310009E030008C",
                INIT_06 => X"0502588FE110E00FE132C04461006001B0000500C005E0006031C005E0016030",
                INIT_07 => X"0501588FE110E00FE132C0446110600F05035886E110E00FE132C0446110600F",
                INIT_08 => X"600F4095E010A000E0FF6010E00F8001E0FF600FE110E00FE132C0446110600F",
                INIT_09 => X"E009600DE008600CE007600B6706E006000006000813E110E00FA13280446110",
                INIT_0A => X"0002A080600C0400C207C106621261118801E01270808801E0117080E00A600E",
                INIT_0B => X"84011400D040000200020002A08060101400D04000020002A080600E1400D040",
                INIT_0C => X"C10662126111E012A000E0FF6012E0118001E0FF601150D12080B01001806010",
                INIT_0D => X"54E34400C401C0050010C005000FE010B01061106012E00F9010610F6011C207",
                INIT_0E => X"0157014F54F14400C40141110174016B0157014754EB4400C401411101740157",
                INIT_0F => X"C4014111016B015754FF4400C4014111016B0157014F014754F94400C4014111",
                INIT_10 => X"0157014F014741110174016B0157014F550D4400C40141110157014755054400",
                INIT_11 => X"E00DB130902063086207610E600DE10CE00BB1309020630A6209610C600B0174",
                INIT_12 => X"B050000251464000B05000034099412A552956F06F2F8601E00680016006E10E",
                INIT_13 => X"E0FF600D51464000B0500001E00CA000E0FF600CE00B8001E0FF600B513A4000",
                INIT_14 => X"B000A000E008E0006008E007E0016007B000417DE00EA000E0FF600EE00D8001",
                INIT_15 => X"6007E008000A6008B000C701516A40001070A000E00AE000600AE009E0016009",
                INIT_16 => X"6008E0078001E0FF6007A0004157E00900086009E00A000A600AB000E0070008",
                INIT_17 => X"600CE003600BA000E00AA000E0FF600AE0098001E0FF6009A000E008A000E0FF",
                INIT_18 => X"6004C0016005C0046003C0046002C0026002C0026003E004600EE005600DE002",
                INIT_19 => X"01B7002801001260030001BA0033010362026303A000C0036005C0036004C001",
                INIT_1A => X"C017603BC016603CE03B01B7002801001260030001BA0033010362046305E03C",
                INIT_1B => X"E10054000600070014201530A000B1309020A000F130D02041B3404BC020003F",
                INIT_1C => X"41D255D459D0520041D451CC59D05310A00041BEA7008601F510D40059C75510",
                INIT_1D => X"0000000000000000000000000000000000000000A000040441D5040241D50401",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"3A503A503A500A28F88E2388E222294088888888888888888888888888888888",
               INITP_01 => X"7FD7FFD7FD7FFD7FD62242428242434042A00A0080A061888882029439090A50",
               INITP_02 => X"229090A4242E8A0A281D2924292439090D09090D0D0FD19294029403FFFFD7FD",
               INITP_03 => X"0000000000000000000008CCFDFDB55D500965F888B00C02C0300A2222222222",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
