--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "0900001209010012090100120903001209050012090A00120913001209200F13";
attribute INIT_01 of ram_1024_x_18  : label is "0F4DEF35EF33EF390F00EF3D0F00EF3E0F00EF10CF13A0008F01F9F040150012";
attribute INIT_02 of ram_1024_x_18  : label is "403350304F686F3DEF3EAF00CF036F3EEF3D8F01CF036F3D0B136A100900EF37";
attribute INIT_03 of ram_1024_x_18  : label is "0F01404B503F44010179005A0100623D633EEF086F3EEF096F3D51874F016F3E";
attribute INIT_04 of ram_1024_x_18  : label is "017900B40100623D633E4088CF086F08CF076F09EF086F3EEF096F3DCF04EF24";
attribute INIT_05 of ram_1024_x_18  : label is "6F08CF076F09E009E108013800B40100623D633ECF04EF240F02406250534401";
attribute INIT_06 of ram_1024_x_18  : label is "613E02B40300CF04EF240F034079506A44010179000E0101623D633E4088CF08";
attribute INIT_07 of ram_1024_x_18  : label is "603D613E020E0301CF04EF240F044088CF086F08CF076F09E009E1080138603D";
attribute INIT_08 of ram_1024_x_18  : label is "CC010F0A50914C001C906F3750C359A04088CF086F08CF076F09E009E1080138";
attribute INIT_09 of ram_1024_x_18  : label is "4480A4806408EF3B7F1011B0EF355496CC010F0A50994C001C906F39EF33548E";
attribute INIT_0A of ram_1024_x_18  : label is "E108E009E100D020623B61086009E039904064336039E037D0406435603750B1";
attribute INIT_0B of ram_1024_x_18  : label is "E108E009A1009020623B61086009E039D04064336039E03790406435603740C0";
attribute INIT_0C of ram_1024_x_18  : label is "40D950D04003602440E2E0378001E0FF603740CC50C74002602440888B018901";
attribute INIT_0D of ram_1024_x_18  : label is "8001E0FF603940E250DD4004602440E2E0398001E0FF6039E0378001E0FF6037";
attribute INIT_0E of ram_1024_x_18  : label is "000A000AC002600BE0228028000A000AC001600DE00D6039E00B603740E2E039";
attribute INIT_0F of ram_1024_x_18  : label is "0125104011601730162015101400401BC020003FC0176023C0166022E0238028";
attribute INIT_10 of ram_1024_x_18  : label is "E107012510501170E004E105012510501160E002E103012510401170E000E101";
attribute INIT_11 of ram_1024_x_18  : label is "670701716400650106000700017100006104620503000400650266030700E006";
attribute INIT_12 of ram_1024_x_18  : label is "040803089310512E3020040003000201E43DE33EE23FA0000171040005006606";
attribute INIT_13 of ram_1024_x_18  : label is "54000600070014201530A000F130D020A000643D633E623F10401130552B0206";
attribute INIT_14 of ram_1024_x_18  : label is "5151596756204165514D59635730A000413FA7008601F510D40059485510E100";
attribute INIT_15 of ram_1024_x_18  : label is "0801416B0804416B0801416B0802415D5159595B540041615155595F55104169";
attribute INIT_16 of ram_1024_x_18  : label is "F370F260F150D040A000416B0804416B0801416B0804416B0801416B0804416B";
attribute INIT_17 of ram_1024_x_18  : label is "5585598152004185517D59815310A000B1309020A000B370B260B1509040A000";
attribute INIT_18 of ram_1024_x_18  : label is "000000000000000000000000000000004187A000040441860402418604014183";
attribute INIT_19 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "00A388AC028F700E22B00A3DC038888A3DC02234F49898022A22266F33333330";
attribute INITP_01 of ram_1024_x_18 : label is "C0038889A89A888E43D39090F4E43D35A5024243A5024243420B6D0B6D0DE22B";
attribute INITP_02 of ram_1024_x_18 : label is "F7F6595655B333333333F7F7F7F6D5754025800EA740AAC0300C0002B0AC2B0A";
attribute INITP_03 of ram_1024_x_18 : label is "000000000000000000000000000000000000000000000000000000000000E333";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"0900001209010012090100120903001209050012090A00120913001209200F13",
                INIT_01 => X"0F4DEF35EF33EF390F00EF3D0F00EF3E0F00EF10CF13A0008F01F9F040150012",
                INIT_02 => X"403350304F686F3DEF3EAF00CF036F3EEF3D8F01CF036F3D0B136A100900EF37",
                INIT_03 => X"0F01404B503F44010179005A0100623D633EEF086F3EEF096F3D51874F016F3E",
                INIT_04 => X"017900B40100623D633E4088CF086F08CF076F09EF086F3EEF096F3DCF04EF24",
                INIT_05 => X"6F08CF076F09E009E108013800B40100623D633ECF04EF240F02406250534401",
                INIT_06 => X"613E02B40300CF04EF240F034079506A44010179000E0101623D633E4088CF08",
                INIT_07 => X"603D613E020E0301CF04EF240F044088CF086F08CF076F09E009E1080138603D",
                INIT_08 => X"CC010F0A50914C001C906F3750C359A04088CF086F08CF076F09E009E1080138",
                INIT_09 => X"4480A4806408EF3B7F1011B0EF355496CC010F0A50994C001C906F39EF33548E",
                INIT_0A => X"E108E009E100D020623B61086009E039904064336039E037D0406435603750B1",
                INIT_0B => X"E108E009A1009020623B61086009E039D04064336039E03790406435603740C0",
                INIT_0C => X"40D950D04003602440E2E0378001E0FF603740CC50C74002602440888B018901",
                INIT_0D => X"8001E0FF603940E250DD4004602440E2E0398001E0FF6039E0378001E0FF6037",
                INIT_0E => X"000A000AC002600BE0228028000A000AC001600DE00D6039E00B603740E2E039",
                INIT_0F => X"0125104011601730162015101400401BC020003FC0176023C0166022E0238028",
                INIT_10 => X"E107012510501170E004E105012510501160E002E103012510401170E000E101",
                INIT_11 => X"670701716400650106000700017100006104620503000400650266030700E006",
                INIT_12 => X"040803089310512E3020040003000201E43DE33EE23FA0000171040005006606",
                INIT_13 => X"54000600070014201530A000F130D020A000643D633E623F10401130552B0206",
                INIT_14 => X"5151596756204165514D59635730A000413FA7008601F510D40059485510E100",
                INIT_15 => X"0801416B0804416B0801416B0802415D5159595B540041615155595F55104169",
                INIT_16 => X"F370F260F150D040A000416B0804416B0801416B0804416B0801416B0804416B",
                INIT_17 => X"5585598152004185517D59815310A000B1309020A000B370B260B1509040A000",
                INIT_18 => X"000000000000000000000000000000004187A000040441860402418604014183",
                INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"00A388AC028F700E22B00A3DC038888A3DC02234F49898022A22266F33333330",
               INITP_01 => X"C0038889A89A888E43D39090F4E43D35A5024243A5024243420B6D0B6D0DE22B",
               INITP_02 => X"F7F6595655B333333333F7F7F7F6D5754025800EA740AAC0300C0002B0AC2B0A",
               INITP_03 => X"000000000000000000000000000000000000000000000000000000000000E333",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
