--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A00D5E019001FE01800B6E017003EE01600B1E0150076E014000FE01300C9";
attribute INIT_01 of ram_1024_x_18  : label is "E02200FFE0210001E02000FFE01F0003E01E00FFE01D0007E01C00FAE01B000F";
attribute INIT_02 of ram_1024_x_18  : label is "E02A001FE0290000E028003FE0270000E026007FE0250000E02400FFE0230000";
attribute INIT_03 of ram_1024_x_18  : label is "E0320001E0310000E0300003E02F0000E02E0007E02D0000E02C000FE02B0000";
attribute INIT_04 of ram_1024_x_18  : label is "8001D01001130032EE3D0E00EE3E0E00ED390D00ED3A0D00EC370C9BEC380C74";
attribute INIT_05 of ram_1024_x_18  : label is "0147623D633EEE3EAE04CE036E3EEE3D8E77CE036E3D0B130A0F0900E010000E";
attribute INIT_06 of ram_1024_x_18  : label is "020A50734300139062386137EF086F3EEF096F3D50E459A051984404018A0058";
attribute INIT_07 of ram_1024_x_18  : label is "E236E135547AC3010108020A507E43001390623A6139E234E133546FC3010108";
attribute INIT_08 of ram_1024_x_18  : label is "603754B14380A380A300E3FF63088201E2FF6209EF3B7F108101EF3C7F1011B0";
attribute INIT_09 of ram_1024_x_18  : label is "6534643303000200613A6039E104E005017D0700060065366435030002006138";
attribute INIT_0A of ram_1024_x_18  : label is "E102E003017D07000600653C643B0300020061086009E106E007018207000600";
attribute INIT_0B of ram_1024_x_18  : label is "03000200613A6039E104E00501820700060065366435030002006138603740D4";
attribute INIT_0C of ram_1024_x_18  : label is "018207000600653C643B0300020061086009E106E007017D0700060065346433";
attribute INIT_0D of ram_1024_x_18  : label is "6F03EF396F07EF3A6F06EF376F05EF386F048B018B018901E102E003CF040FFF";
attribute INIT_0E of ram_1024_x_18  : label is "C302C202620B630AE00C603AE00D6039E00A6038E00B60374064EF086F02EF09";
attribute INIT_0F of ram_1024_x_18  : label is "014C00330103C301C201620D630CE03C01870028010012600300014C00330103";
attribute INIT_10 of ram_1024_x_18  : label is "1620151014004052C020003FC017603BC016603CE03B0187002801A912600300";
attribute INIT_11 of ram_1024_x_18  : label is "E004E105013910501160E002E103013910401170E000E1010139104011601730";
attribute INIT_12 of ram_1024_x_18  : label is "06000700018200006104620503000400650266030700E006E107013910501170";
attribute INIT_13 of ram_1024_x_18  : label is "3020040003000201E43DE33EE23FA00001820400050066066707018264006501";
attribute INIT_14 of ram_1024_x_18  : label is "0600070014201530A000643D633E623F10401130553F02060408030893105142";
attribute INIT_15 of ram_1024_x_18  : label is "597856204176515E59745730A0004150A7008601F510D40059595510E1005400";
attribute INIT_16 of ram_1024_x_18  : label is "417C0804417C0801417C0802416E516A596C54004172516659705510417A5162";
attribute INIT_17 of ram_1024_x_18  : label is "F260F150D040A000417C0804417C0801417C0804417C0801417C0804417C0801";
attribute INIT_18 of ram_1024_x_18  : label is "599252004196518E59925310A000B1309020A000B370B260B1509040A000F370";
attribute INIT_19 of ram_1024_x_18  : label is "00000000000000000000000000004198A0000404419704024197040141945596";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "ADAD02B6B4088DDC0262600A5088888888888888888888888888888888888888";
attribute INITP_01 of ram_1024_x_18 : label is "C282C030A08888E2222215A8C0002B0000AC0003AC0002B0000AC00034410860";
attribute INITP_02 of ram_1024_x_18 : label is "56CCCCCCCCCFDFDFDFDB55D500800EA740AAC0300C0002B0AC2B0AC003888B00";
attribute INITP_03 of ram_1024_x_18 : label is "00000000000000000000000000000000000000000000000000038CCFDFD96559";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A00D5E019001FE01800B6E017003EE01600B1E0150076E014000FE01300C9",
                INIT_01 => X"E02200FFE0210001E02000FFE01F0003E01E00FFE01D0007E01C00FAE01B000F",
                INIT_02 => X"E02A001FE0290000E028003FE0270000E026007FE0250000E02400FFE0230000",
                INIT_03 => X"E0320001E0310000E0300003E02F0000E02E0007E02D0000E02C000FE02B0000",
                INIT_04 => X"8001D01001130032EE3D0E00EE3E0E00ED390D00ED3A0D00EC370C9BEC380C74",
                INIT_05 => X"0147623D633EEE3EAE04CE036E3EEE3D8E77CE036E3D0B130A0F0900E010000E",
                INIT_06 => X"020A50734300139062386137EF086F3EEF096F3D50E459A051984404018A0058",
                INIT_07 => X"E236E135547AC3010108020A507E43001390623A6139E234E133546FC3010108",
                INIT_08 => X"603754B14380A380A300E3FF63088201E2FF6209EF3B7F108101EF3C7F1011B0",
                INIT_09 => X"6534643303000200613A6039E104E005017D0700060065366435030002006138",
                INIT_0A => X"E102E003017D07000600653C643B0300020061086009E106E007018207000600",
                INIT_0B => X"03000200613A6039E104E00501820700060065366435030002006138603740D4",
                INIT_0C => X"018207000600653C643B0300020061086009E106E007017D0700060065346433",
                INIT_0D => X"6F03EF396F07EF3A6F06EF376F05EF386F048B018B018901E102E003CF040FFF",
                INIT_0E => X"C302C202620B630AE00C603AE00D6039E00A6038E00B60374064EF086F02EF09",
                INIT_0F => X"014C00330103C301C201620D630CE03C01870028010012600300014C00330103",
                INIT_10 => X"1620151014004052C020003FC017603BC016603CE03B0187002801A912600300",
                INIT_11 => X"E004E105013910501160E002E103013910401170E000E1010139104011601730",
                INIT_12 => X"06000700018200006104620503000400650266030700E006E107013910501170",
                INIT_13 => X"3020040003000201E43DE33EE23FA00001820400050066066707018264006501",
                INIT_14 => X"0600070014201530A000643D633E623F10401130553F02060408030893105142",
                INIT_15 => X"597856204176515E59745730A0004150A7008601F510D40059595510E1005400",
                INIT_16 => X"417C0804417C0801417C0802416E516A596C54004172516659705510417A5162",
                INIT_17 => X"F260F150D040A000417C0804417C0801417C0804417C0801417C0804417C0801",
                INIT_18 => X"599252004196518E59925310A000B1309020A000B370B260B1509040A000F370",
                INIT_19 => X"00000000000000000000000000004198A0000404419704024197040141945596",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"ADAD02B6B4088DDC0262600A5088888888888888888888888888888888888888",
               INITP_01 => X"C282C030A08888E2222215A8C0002B0000AC0003AC0002B0000AC00034410860",
               INITP_02 => X"56CCCCCCCCCFDFDFDFDB55D500800EA740AAC0300C0002B0AC2B0AC003888B00",
               INITP_03 => X"00000000000000000000000000000000000000000000000000038CCFDFD96559",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
