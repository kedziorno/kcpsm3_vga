--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E01A0000E0190001E0180001E0170003E0160005E015000AE0140013E0130020";
attribute INIT_01 of ram_1024_x_18  : label is "0A080900ED390D00EC370C4DE010000E8001D0100113001AEE3D0E00EE3E0E00";
attribute INIT_02 of ram_1024_x_18  : label is "0100623D633EEF086F3EEF096F3DEE3EAE00CE036E3EEE3D8E01CE036E3D0B13";
attribute INIT_03 of ram_1024_x_18  : label is "0100623D633E406EEF086F3EEF096F3DC004E0240001403D503544010156005A";
attribute INIT_04 of ram_1024_x_18  : label is "406EE009E1080115603D613E02B40300C004E0240002405050454401015600B4";
attribute INIT_05 of ram_1024_x_18  : label is "011500B40100023D033EC004E02400034063505844010156000E0101623D633E";
attribute INIT_06 of ram_1024_x_18  : label is "50A959A0E208A200E2FF623EE2098201E2FF623DC004E0240004406EE009E108";
attribute INIT_07 of ram_1024_x_18  : label is "E135547CC301010A507F430013906139E1335474C301010A5077430013906137";
attribute INIT_08 of ram_1024_x_18  : label is "6009E039904064336039E037D0406435603750974480A4806408EF3B7F1011B0";
attribute INIT_09 of ram_1024_x_18  : label is "6009E039D04064336039E03790406435603740A6E108E009E100D020623B6108";
attribute INIT_0A of ram_1024_x_18  : label is "603740B450AF400450AF40016024406E8B018901E108E009A1009020623B6108";
attribute INIT_0B of ram_1024_x_18  : label is "603740BFE0398001E0FF603940BF50BA400250BA4001602440BFE0378001E0FF";
attribute INIT_0C of ram_1024_x_18  : label is "6022E0238028000A000AC002600BE0228028000A000AC001600DE00D6039E00B";
attribute INIT_0D of ram_1024_x_18  : label is "1170E000E1010102104011601730162015101400401AC020003FC0176023C016";
attribute INIT_0E of ram_1024_x_18  : label is "66030700E006E107010210501170E004E105010210501160E002E10301021040";
attribute INIT_0F of ram_1024_x_18  : label is "0400050066066707014E6400650106000700014E000061046205030004006502";
attribute INIT_10 of ram_1024_x_18  : label is "113055080206040803089310510B3020040003000201E43DE33EE23FA000014E";
attribute INIT_11 of ram_1024_x_18  : label is "59255510E10054000600070014201530A000F130D020A000643D633E623F1040";
attribute INIT_12 of ram_1024_x_18  : label is "593C55104146512E594456204142512A59405730A000411CA7008601F510D400";
attribute INIT_13 of ram_1024_x_18  : label is "4148080441480801414808044148080141480802413A513659385400413E5132";
attribute INIT_14 of ram_1024_x_18  : label is "B1509040A000F370F260F150D040A00041480804414808014148080441480801";
attribute INIT_15 of ram_1024_x_18  : label is "4163040141605562595E52004162515A595E5310A000B1309020A000B370B260";
attribute INIT_16 of ram_1024_x_18  : label is "000000000000000000000000000000000000000000004164A000040441630402";
attribute INIT_17 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_18 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_19 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "B6D0B6D0D9090A3AC028F700EB00A3DC0388A3DC02226260088A508888888888";
attribute INITP_01 of ram_1024_x_18 : label is "00C030000AC2B0AC2B000E2226A26A22390F74E43DD35A5024243A5024243420";
attribute INITP_02 of ram_1024_x_18 : label is "000000000000038CCFDFD9655956CCCCCCCCCFDFDFDFDB55D50096003A9D02AB";
attribute INITP_03 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E01A0000E0190001E0180001E0170003E0160005E015000AE0140013E0130020",
                INIT_01 => X"0A080900ED390D00EC370C4DE010000E8001D0100113001AEE3D0E00EE3E0E00",
                INIT_02 => X"0100623D633EEF086F3EEF096F3DEE3EAE00CE036E3EEE3D8E01CE036E3D0B13",
                INIT_03 => X"0100623D633E406EEF086F3EEF096F3DC004E0240001403D503544010156005A",
                INIT_04 => X"406EE009E1080115603D613E02B40300C004E0240002405050454401015600B4",
                INIT_05 => X"011500B40100023D033EC004E02400034063505844010156000E0101623D633E",
                INIT_06 => X"50A959A0E208A200E2FF623EE2098201E2FF623DC004E0240004406EE009E108",
                INIT_07 => X"E135547CC301010A507F430013906139E1335474C301010A5077430013906137",
                INIT_08 => X"6009E039904064336039E037D0406435603750974480A4806408EF3B7F1011B0",
                INIT_09 => X"6009E039D04064336039E03790406435603740A6E108E009E100D020623B6108",
                INIT_0A => X"603740B450AF400450AF40016024406E8B018901E108E009A1009020623B6108",
                INIT_0B => X"603740BFE0398001E0FF603940BF50BA400250BA4001602440BFE0378001E0FF",
                INIT_0C => X"6022E0238028000A000AC002600BE0228028000A000AC001600DE00D6039E00B",
                INIT_0D => X"1170E000E1010102104011601730162015101400401AC020003FC0176023C016",
                INIT_0E => X"66030700E006E107010210501170E004E105010210501160E002E10301021040",
                INIT_0F => X"0400050066066707014E6400650106000700014E000061046205030004006502",
                INIT_10 => X"113055080206040803089310510B3020040003000201E43DE33EE23FA000014E",
                INIT_11 => X"59255510E10054000600070014201530A000F130D020A000643D633E623F1040",
                INIT_12 => X"593C55104146512E594456204142512A59405730A000411CA7008601F510D400",
                INIT_13 => X"4148080441480801414808044148080141480802413A513659385400413E5132",
                INIT_14 => X"B1509040A000F370F260F150D040A00041480804414808014148080441480801",
                INIT_15 => X"4163040141605562595E52004162515A595E5310A000B1309020A000B370B260",
                INIT_16 => X"000000000000000000000000000000000000000000004164A000040441630402",
                INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"B6D0B6D0D9090A3AC028F700EB00A3DC0388A3DC02226260088A508888888888",
               INITP_01 => X"00C030000AC2B0AC2B000E2226A26A22390F74E43DD35A5024243A5024243420",
               INITP_02 => X"000000000000038CCFDFD9655956CCCCCCCCCFDFDFDFDB55D50096003A9D02AB",
               INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
