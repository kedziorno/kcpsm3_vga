--
-- Definition of a single port ROM for KCPSM3 program defined by program.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity program is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end program;
--
architecture low_level_definition of program is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E7070709E706070EE7050790E704071AE7030700E702072DE701079BE7000700";
attribute INIT_01 of ram_1024_x_18  : label is "E70F07E5E70E0700E70D07CBE70C0701E70B0793E70A0703E7090720E7080707";
attribute INIT_02 of ram_1024_x_18  : label is "CE03CD03AF00AE008DFF0D000E000F00E713073AE7120700E7110772E7100700";
attribute INIT_03 of ram_1024_x_18  : label is "0700C7040701C1064801013910D011E012F003000400056806010700C105CF03";
attribute INIT_04 of ram_1024_x_18  : label is "070216F015E014D0E739070150514804013910D011E012F00300040005010600";
attribute INIT_05 of ram_1024_x_18  : label is "06000700E7390702506C4804013910D011E012F003000400050206000700C704";
attribute INIT_06 of ram_1024_x_18  : label is "0400050306000700C704070316F015E014D0015C10D011E012F0030004000502";
attribute INIT_07 of ram_1024_x_18  : label is "01020200030014D015E016F00700E739070350874804013910D011E012F00300";
attribute INIT_08 of ram_1024_x_18  : label is "A700E7FF17E01D708701E7FF17D0E7390704C704070416F015E014D0015C0000";
attribute INIT_09 of ram_1024_x_18  : label is "E73807FF708088017180080016F015E014D0C70407051F70A700E7FF17F01E70";
attribute INIT_0A of ram_1024_x_18  : label is "0A08090A50B4470067381C201B301A001910E73887016738C7040707C7040706";
attribute INIT_0B of ram_1024_x_18  : label is "79808801B39092A0F1B0D0C054C8A780176050E04709673840ACC7010C080B0A";
attribute INIT_0C of ram_1024_x_18  : label is "7A80880179808801F390D2A0B1B090C040A2C70407EEE600F590D4A07A808801";
attribute INIT_0D of ram_1024_x_18  : label is "40E0020003010000010040E0020003000000010140A2C70407FFA600B59094A0";
attribute INIT_0E of ram_1024_x_18  : label is "673940FE1170A700E7FF171010708701E7FF170040EF50E6470450E647016739";
attribute INIT_0F of ram_1024_x_18  : label is "E13EE03F40FE1370A700E7FF173012708701E7FF172040FE50F5470250F54701";
attribute INIT_10 of ram_1024_x_18  : label is "0A08090A0A08090A0A08090A0A08090A0A08090AC902CA026A3F693EE33CE23D";
attribute INIT_11 of ram_1024_x_18  : label is "8A280A08090A0A08090A0A08090A0A08090A0A08090AC901CA016A3D693CEA3B";
attribute INIT_12 of ram_1024_x_18  : label is "52700400080012001530A000B1309700402BC720073FC717673AC716673BEA3A";
attribute INIT_13 of ram_1024_x_18  : label is "5141595756204155513D59535730A000412FA8008401F510D27059385510E100";
attribute INIT_14 of ram_1024_x_18  : label is "0801415B0804415B0801415B0802414D5149594B540041515145594F55104159";
attribute INIT_15 of ram_1024_x_18  : label is "F370F260F150D040A000415B0804415B0801415B0804415B0801415B0804415B";
attribute INIT_16 of ram_1024_x_18  : label is "000000000000000000000000000000000000000000000000000000004161A000";
attribute INIT_17 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_18 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_19 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "000237000080300008DC0002008DC0002270000AA54088888888888888888888";
attribute INITP_01 of ram_1024_x_18 : label is "AC4043DD31010F74C0300E151155E151155C34DAAD002488810020404042200C";
attribute INITP_02 of ram_1024_x_18 : label is "000000000000000E55B333333333F7F7F7F6D5754025E2226AAAAA82AAAAAA0A";
attribute INITP_03 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E7070709E706070EE7050790E704071AE7030700E702072DE701079BE7000700",
                INIT_01 => X"E70F07E5E70E0700E70D07CBE70C0701E70B0793E70A0703E7090720E7080707",
                INIT_02 => X"CE03CD03AF00AE008DFF0D000E000F00E713073AE7120700E7110772E7100700",
                INIT_03 => X"0700C7040701C1064801013910D011E012F003000400056806010700C105CF03",
                INIT_04 => X"070216F015E014D0E739070150514804013910D011E012F00300040005010600",
                INIT_05 => X"06000700E7390702506C4804013910D011E012F003000400050206000700C704",
                INIT_06 => X"0400050306000700C704070316F015E014D0015C10D011E012F0030004000502",
                INIT_07 => X"01020200030014D015E016F00700E739070350874804013910D011E012F00300",
                INIT_08 => X"A700E7FF17E01D708701E7FF17D0E7390704C704070416F015E014D0015C0000",
                INIT_09 => X"E73807FF708088017180080016F015E014D0C70407051F70A700E7FF17F01E70",
                INIT_0A => X"0A08090A50B4470067381C201B301A001910E73887016738C7040707C7040706",
                INIT_0B => X"79808801B39092A0F1B0D0C054C8A780176050E04709673840ACC7010C080B0A",
                INIT_0C => X"7A80880179808801F390D2A0B1B090C040A2C70407EEE600F590D4A07A808801",
                INIT_0D => X"40E0020003010000010040E0020003000000010140A2C70407FFA600B59094A0",
                INIT_0E => X"673940FE1170A700E7FF171010708701E7FF170040EF50E6470450E647016739",
                INIT_0F => X"E13EE03F40FE1370A700E7FF173012708701E7FF172040FE50F5470250F54701",
                INIT_10 => X"0A08090A0A08090A0A08090A0A08090A0A08090AC902CA026A3F693EE33CE23D",
                INIT_11 => X"8A280A08090A0A08090A0A08090A0A08090A0A08090AC901CA016A3D693CEA3B",
                INIT_12 => X"52700400080012001530A000B1309700402BC720073FC717673AC716673BEA3A",
                INIT_13 => X"5141595756204155513D59535730A000412FA8008401F510D27059385510E100",
                INIT_14 => X"0801415B0804415B0801415B0802414D5149594B540041515145594F55104159",
                INIT_15 => X"F370F260F150D040A000415B0804415B0801415B0804415B0801415B0804415B",
                INIT_16 => X"000000000000000000000000000000000000000000000000000000004161A000",
                INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"000237000080300008DC0002008DC0002270000AA54088888888888888888888",
               INITP_01 => X"AC4043DD31010F74C0300E151155E151155C34DAAD002488810020404042200C",
               INITP_02 => X"000000000000000E55B333333333F7F7F7F6D5754025E2226AAAAA82AAAAAA0A",
               INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE program.vhd
--
------------------------------------------------------------------------------------
